-- EECS 361 Pipelined Processor
-- This calculates the inputs to be fed into the EX stage



