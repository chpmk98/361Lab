-- EECS 361 Single-Cycle Processor
-- by Alvin Tan

-- An unfortunate series of huge muxes necessary to determine which register is outputted to 
-- busA and busB in reg_comp.
-- Input: 32 32-bit values

entity reg_32to1mux is
end reg_32to1mux;






